module BCD_DECO(N, a, b, c, d, e, f, g);
    input N[3:0];
    output a, b, c, d, e, f, g;

    always @(N) begin

    end

endmodule