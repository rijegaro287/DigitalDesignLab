module unidad_logica();

endmodule