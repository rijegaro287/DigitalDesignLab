module unidad_arimetica();

endmodule