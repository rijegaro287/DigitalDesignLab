module instruction_memory(
  input logic [31:0] addr,
  output logic [31:0] data
);

endmodule

// 11100101100100000000000000000000; // LDR R0, [R0], #0x00
// b11100101100100010001000000000001; // LDR R1, [R1], #0x01
// b11100101100100000010000000000010; // LDR R2, [R0], #0x02

// 1110 00 1 0100 0 0000 0000 0000 00000010 // ADD R0, R0, #0x02
// 1110 00 1 0100 0 0000 0001 0000 00000101 // ADD R1, R0, #0x05
// 1110 00 1 0100 0 0001 0010 0000 00101010 // ADD R2, R1, #0x2A
// 1110 00 0 0100 0 0010 0001 00000 00 0 0000 // ADD R1, R2, R0
// 1110 00 0 0100 0 0010 0010 00000 00 0 0010 // ADD R2, R2, R2