module datapath_tb();

endmodule