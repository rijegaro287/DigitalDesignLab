module main(
  input logic clk,
  input logic rst
);

endmodule