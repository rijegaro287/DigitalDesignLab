module BCD_DECO_TB();
    reg N[3:0];
    wire a, b, c, d, e, f, g;


endmodule