module BCD_DECO_TB();
    reg N[3:0];
    wire BCD[6:0];


endmodule